library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity x_cor is
  port(rst_n: in std_logic;
       clk: in std_logic;
       din: in std_logic_vector(11 downto 0);
       dout1:out std_logic_vector(20 downto 0);
       dout2:out std_logic_vector(20 downto 0));
end entity x_cor;

architecture rtl of x_cor is
   --signal tmp: std_logic_vector(11 downto 0);
   --signal tmp1: std_logic_vector(19 downto 0);
   component reg_12 is
   port(rst_n: in std_logic;
        clk: in std_logic;
        din: in std_logic_vector(11 downto 0);
        do:out std_logic_vector(11 downto 0));
end component reg_12;
type ram is array (0 to 255) of std_logic_vector(11 downto 0);--255
signal reg,reg1,reg2: ram;
type ram1 is array (0 to 255) of std_logic_vector(20 downto 0);--255
signal reg3,reg4:ram1;
type rom is array (255 downto 0) of std_logic; --255
--constant coef: rom:=( '1','1','1','1','0','0','0','0','1','1','1','1','1','1','0','0',
--                      '0','0','0','1','1','1','1','1','0','0','0','0','0','1','1','1',
--                      '1','1','0','0','0','0','1','1','1','1','1','0','0','0','0','1',	
--                      '1','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0');
--constant coef: rom:=(  '1','1','1','1','1','1','1','1','0','0','0','0','0','0','1','1',
--							  '1','1','0','0','0','1','1','1','0','0','1','1','0','0','1','1',
--							  '0','0','1','1','0','1','1','0','1','1','0','1','1','0','1','0',
--							  '1','1','0','1','0','1','0','1','1','1','1','1','1','1','1','1');
--constant coef: rom:=('1','1','1','1','1','1','1','1','1','0','0','0','0','0','1','1',	
--                     '1','1','0','0','0','1','1','0','0','0','1','1','0','0','1','1',	
--							'1','0','0','1','1','1','0','1','1','1','0','0','1','1','1','1',	
--							'1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1'); 
--constant coef: rom:=('1','1','1','0','0','0','1','1','1','0','0','0','1','1','0','0',
--                   	'1','1','0','0','1','1','0','1','1','0','1','1','0','0','1','0',	
--							'0','1','1','0','1','0','0','1','0','0','1','0','0','1','1','0',	
--							'1','0','0','0','0','1','1','1','1','1','0','0','0','0','0','1');--for M=8					
--constant coef: rom:=('1','1','0','0','1','1','1','0','0','1','1','0','0','1','1','0',	
--                     '1','1','0','1','1','0','1','1','0','1','0','1','1','0','1','0',	
--							'0','1','0','1','0','0','1','0','1','1','0','1','0','1','1','1',	
--							'1','0','0','1','1','1','0','0','0','0','1','1','1','0','0','1');	--FOR M=12		
--constant coef: rom:=('1','1','0','0','1','1','0','0','1','1','0','0','1','0','1','1',	
--                     '0','0','1','0','0','1','0','0','1','0','0','1','0','1','1','0',	
--							'0','1','0','1','0','0','1','1','0','1','0','0','1','0','0','0',	
--							'0','1','1','0','0','1','1','1','0','0','1','1','1','1','0','0');	--for M=14,10 CARRIERS		
			
constant coef: rom:=('1','1','1','1','0','0','1','1','1','1','1','0','0','0','1','1',
                   	'1','1','0','0','0','1','1','1','1','0','0','0','0','1','1','1',	
							'0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0',	
							'0','1','1','1','1','0','0','0','1','1','1','0','0','0','1','1',	
							'1','0','0','0','0','1','1','1','0','0','0','1','1','1','0','0',
							'0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','1',	
							'0','0','1','1','1','0','0','0','1','1','1','0','0','1','1','1',	
							'0','0','0','1','1','1','0','0','1','1','1','0','0','1','1','1',
							'0','0','0','1','1','0','0','0','1','1','0','0','0','1','1','0',	
							'0','0','1','1','0','0','0','1','1','0','0','0','1','1','0','0',
							'1','1','1','0','0','1','1','1','0','0','1','1','0','0','1','1',	
							'1','0','0','1','1','0','0','1','1','1','0','0','1','1','0','0',	
							'1','1','1','0','0','1','1','0','0','1','1','0','0','0','1','1',	
							'0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','1',	
							'1','0','1','1','0','0','0','1','1','0','0','1','0','0','0','1',	
							'1','0','1','1','0','0','0','1','1','0','1','1','0','0','0','1');--for M=23,C=36 
 
 begin
  reg(0)<=din;
  g1: for i in 0 to 254 generate --254
      u1: reg_12 port map(rst_n,clk,reg(i),reg(i+1));   
  end generate;
      process(reg)is
       begin
             for i in 0 to 255 loop --255
                if coef(i)='0' then
							reg1(i)<=0-reg(i);
                else
                    reg1(i)<=reg(i);
                end if;
					 reg3(i)<=reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i)(11)&reg1(i);
              end loop;
        end process;
        
        process(rst_n,clk) is
          variable tmp: std_logic_vector(20 downto 0);
          begin
			 if rst_n='0' then
			   dout1<=(others=>'0');
          elsif clk'event and clk='1' then
            tmp:=(others=>'0');
            for i in 0 to 255 loop --255
             tmp:=tmp+reg3(i);
            end loop;
            dout1<=tmp;
          end if;
        end process;  

       
 
      process(reg)is
       begin
             for i in 0 to 255 loop --255
                if reg(i)(11)='1' then
                     reg2(i)<=0-reg(i);
                else
                     reg2(i)<=reg(i);
                end if;
					 reg4(i)<=reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i)(11)&reg2(i);
              end loop;
        end process;  
      
      process(rst_n,clk) is
          variable tmp: std_logic_vector(20 downto 0);
          begin
			 if rst_n='0' then
			  dout2<=(others=>'0');
          elsif clk'event and clk='1' then
            tmp:=(others=>'0');
            for i in 0 to 255 loop --255
             tmp:=tmp+reg4(i);
            end loop;
            dout2<=tmp;
          end if;
        end process;  
                 
end architecture rtl;
         
       